`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:51:56 11/30/2016 
// Design Name: 
// Module Name:    Main 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Main();
//-------------------------------------------Entradas-----------------------------------------//
//--------------------------------------------Salidas-----------------------------------------//
//---------------------------------------------Wires------------------------------------------//
	/*wire Read_Data_OutputMEM_to_Read_Data_InputLATCH_MEMWB;
	wire ALU_Result_OutputLATCH_EXMEM_to_ALU_Result_InputLATCH_MEMWB;
	wire Read_Data_OutputLATCH_MEMWB_to_Dato1_InputWB;
	wire ALU_Result_OutputLATCH_MEMWB_to_Dato0_InputWB;*/
//-------------------------------------------Registros----------------------------------------//
//-----------------------------------------Inicializacion-------------------------------------//
//--------------------------------------Declaracion de Bloques--------------------------------//
	/*Main_IF main_if();

	Latch_IF_ID latch_if_id();

	Main_ID main_id();

	Latch_ID_EX latch_id_ex();

	Main_EX main_ex();

	Latch_EX_MEM latch_ex_mem();

	Main_MEM main_mem();

	Latch_MEM_WB latch_mem_wb( Read_Data_OutputMEM_to_Read_Data_InputLATCH_MEMWB,
										ALU_Result_OutputLATCH_EXMEM_to_ALU_Result_InputLATCH_MEMWB,
										Read_Data_OutputLATCH_MEMWB_to_Dato1_InputWB,
										ALU_Result_OutputLATCH_MEMWB_to_Dato0_InputWB );

	Main_WB main_wb(  Read_Data_OutputLATCH_MEMWB_to_Dato1_InputWB,
							ALU_Result_OutputLATCH_MEMWB_to_Dato0_InputWB );*/
//--------------------------------------------Logica------------------------------------------//
endmodule
