`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    00:20:24 12/03/2016 
// Design Name: 
// Module Name:    Instruction_Memory 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Instruction_Memory(addr, read_data);
//-------------------------------------------Entradas-----------------------------------------//
	input [5:0] addr;
//--------------------------------------------Salidas-----------------------------------------//
	output [31:0] read_data;
//---------------------------------------------Wires------------------------------------------//
//-------------------------------------------Registros----------------------------------------//
	reg [31:0] RAM[63:0];
//-----------------------------------------Inicializacion-------------------------------------//
	initial
		begin
			$readmemh("memfile.dat", RAM);
		end
//--------------------------------------Declaracion de Bloques--------------------------------//
//--------------------------------------------Logica------------------------------------------//
	assign read_data = RAM[addr];
endmodule
